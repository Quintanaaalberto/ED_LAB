library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all; -- for addition & counting
use ieee.numeric_std.all;        -- for type conversions

entity Sumador_Restador5Bits is
	port (
		a, b 	: in std_logic_vector(4 downto 0);
		s 		: out std_logic_vector(4 downto 0);
		c_out 	: out std_logic;
		s_r : in std_logic
	) ;
end Sumador_Restador5Bits;

architecture Sumador_Restador5Bits_arc of Sumador_Restador5Bits is
-- intermidiate carries are stored on this vector
	signal c 	: std_logic_vector (5 downto 0);
-- generation and spread, g and p
	signal g, p : std_logic_vector (4 downto 0);
	signal b_j : std_logic_vector(4 downto 0);
	

-- now we reference the other blocks used on the hierarchy
	component Sumador1Bit
	port (
		a_i , b_i 	: in std_logic;
		c_i 		: in std_logic;
		s_i 		: out std_logic;
		p_i , g_i 	: out std_logic);
	end component;

	component CarryLookAhead
	port(
		g, p 		: in std_logic_vector(4 downto 0);
		c_0 		: in std_logic;
		c 			: out std_logic_vector(5 downto 1));
	end component;

begin
	
	process(s_r)
	
		begin 
			if s_r = '0' then 
				c(0) <= '0';
			else 
				c(0) <= '1';
			end if;
	end process;
	
	c_out <= c(5) xor c(4);

	GenSum : for i in 0 to 4 generate
	
		b_j(i) <= b(i) xor s_r;
		
		i_Sumador1Bit : Sumador1Bit
		port map (
			a_i => a(i),
			b_i => b_j(i),
			c_i => c(i),
			s_i => s(i),
			p_i => p(i),
			g_i => g(i)
			);
	end generate GenSum;
-- instanciamos con los vectores de g y p una 
-- ejecución de la operación Carry Look Ahead
	i_CarryLookAhead : CarryLookAhead
	port map (
		g => g,
		p => p,
		c_0 => c(0),
		c => c(5 downto 1));


end  Sumador_Restador5Bits_arc;