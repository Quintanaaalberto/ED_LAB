library ieee;
use ieee.numeric_std.all;
use ieee.std_logic_1164.all;

entity Pr10 is 
	port(
		
		)